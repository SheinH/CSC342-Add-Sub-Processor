    Mac OS X            	   2   q      �                                      ATTR       �   �                     �     com.apple.provenance  s��wu��